//%%%%%%%%%%%%%%%%%%%%%%%%%%%%ALU Test Module%%%%%%%%%%%%%%%%%%%%%%%%
//********************************************************************
//-------------------------------------------------------------------


module ALU_Test_V1;

//local variables
//--------------input
reg [31:0] A,B; 		//32 bit input operands
reg [3:0] OP; 			//Input operation 
reg	CIN; 				//input carry
//--------------output
wire[31:0] R; 			//32-bit ALU result
wire  C,V,N,Z;			//condition codes


//-----------------ARM Instruction set definition---------------------

	parameter  AND = 4'b0000;
	parameter  EOR = 4'b0001;
	parameter  SUB = 4'b0010;
	parameter  RSB = 4'b0011;
	parameter  ADD = 4'b0100;
	parameter  ADC = 4'b0101;
	parameter  SBC = 4'b0110;
	parameter  RSC = 4'b0111;
	parameter  TST = 4'b1000;
	parameter  CMP = 4'b1010;
	parameter  CMN = 4'b1011;
	parameter  ORR = 4'b1100;
	parameter  TEQ = 4'b1001;
	parameter  MOV = 4'b1101;
	parameter  BIC = 4'b1110;
	parameter  MVN = 4'b1111;




//simulation parameters
parameter sim_time = 100000;	//simulation time

ALU_V1 ALU(R,C,Z,V,N,A,B,CIN,OP);		//ALU module instantiation
initial #sim_time $finish;		//simulation termination time

initial	begin
	//initializing inputs
	CIN = 0;		//Input Carry equals 0
	A = 0; B = 0;
	//--------------------------------AND	
	OP = AND;			
	#10; A = 32'h12344567; B = 32'h0000FE18;
	#10; A = 32'h005AC023; B = 32'h0DAE2310;
	#10;
	$display("**********************************************************************");
	//--------------------------------EOR
	OP = EOR; 
	#10; A = 32'h000F000F; B = 32'hFFFFAAFA;
	#10; A = 32'h12344567; B = 32'h0000FE18;

	#10;
	$display("**********************************************************************");
	//--------------------------------SUB
	OP = SUB; 
	#10; A = 32'h005AC023; B = 32'h0DAE2310;
	#10; A = 32'h50000000; B = 32'hB0000000;
	#10;
	$display("**********************************************************************");
	//--------------------------------RSB
	OP = RSB; 
	#10; A = 32'h12344567; B = 32'hF000FE18;
	#10; A = 32'h005AC023; B = 32'h0DAE2310;

	#10;
	$display("**********************************************************************");
	//--------------------------------ADD
	OP = ADD; 
	#10; A = 32'h12344567; B = 32'hF000FE18;
	#10; A = 32'h7F000000; B = 32'h0F001000;  //testing V
	#10;
	$display("**********************************************************************");
	//--------------------------------TST
	OP = TST; 
	#10; A = 32'h12344567; B = 32'h0000FE18;
	#10; A = 32'h005AC023; B = 32'h0DAE2310;

	#10;
	$display("**********************************************************************");
	//--------------------------------TEQ
	OP = TEQ; 
	#10; A = 32'h12344567; B = 32'h0000FE18;
	
	#10;
	$display("**********************************************************************");
	//--------------------------------CMP
	OP = CMP; 
	#10; A = 32'h50000000; B = 32'hB0000000;
	#10;
	$display("**********************************************************************");
	//--------------------------------CMN
	OP = CMN; 
	#10; A = 32'h12344567; B = 32'h0000FE18;
	#10; A = 32'h005AC023; B = 32'h0DAE2310;

	#10;
	$display("**********************************************************************");
	//--------------------------------ORR
	OP = ORR; 
	#10; A = 32'h12344567; B = 32'h0000FE18;

	#10;
	$display("**********************************************************************");
	//--------------------------------MOV
	OP = MOV; 
	#10; A = 32'h005AC023; B = 32'h0DAE2310;

	#10;
	$display("**********************************************************************");
	//--------------------------------BIC
	OP = BIC; 
	#10; A = 32'h12344567; B = 32'h0000FE18;

	#10;
	$display("**********************************************************************");
	//--------------------------------MVN
	OP = MVN; 
	#10; A = 32'h005AC023; B = 32'h0DAE2310;
	#10;

	//-----------------------------------Operation involving Carry bit
	CIN=0;
		$display("**********************************************************************");
		//--------------------------------ADC
		OP = ADC; 
		#10; A = 32'h12344567; B = 32'hF000FE18;
		#10;

		$display("**********************************************************************");
		//--------------------------------SBC
		OP = SBC; 
		#10; A = 32'h005AC023; B = 32'h0DAE2310;
		#10; A = 32'h50000000; B = 32'hB0000000;
		#10;

		$display("**********************************************************************");
		//--------------------------------RSC
		OP = RSC; 
		#10; A = 32'h12344567; B = 32'hF000FE18;
		#10;

	CIN = 1;
		$display("**********************************************************************");
		//--------------------------------ADC
		OP = ADC; 
		#10; A = 32'h50000000; B = 32'hB0000000;
		#10; A = 32'h005AC023; B = 32'h0DAE2310;
		#10;

		$display("**********************************************************************");
		//--------------------------------SBC
		OP = SBC; 
		#10; A = 32'h12344567; B = 32'hF000FE18;
		#10; A = 32'h50000000; B = 32'hB0000000;
		#10;

		$display("**********************************************************************");
		//--------------------------------RSC
		OP = RSC; 
		#10; A = 32'h12344567; B = 32'hF000FE18;
		#10; A = 32'h005AC023; B = 32'h0DAE2310;
		#10;		






end

initial begin 
	$display(" OP   A        B        CIN Result   Z N V C 	   	      Time");		//prints header
	$display("**********************************************************************");
	$monitor(" %b %h %h %b   %h %b %b %b %b %d", OP, A, B, CIN, R, Z, N, V, C, $time);		//print signals
end

endmodule

