
//---------------------ROM 2^8 cells of 64 bits----------------------
module rom (output reg [63:0] OUT, input [7:0] IN);
	
	//IN contains a codified instruction
	//OUT will provde an array of all control variables needed to execute an instruction
	//The format is the following:
	
	//63     62   61   60   59   58     57     56-54   53  52  51  50-48  47    46     45    44      43    42   41  40   39   38   37   36   35   34   33   32   31   30   29  28   27  26   25   24   23      22        21       20    19   18     17      16      15-8      7-0
	//                                         N2-N0  INV  MS  MI  S2-S0  FRLd  RFLd  IRLd  MARLd  MDRLd  R/W  MOV  DS1  DS0  CIN  MA1  MA0  MB2  MB1  MB0  MC2  MC1  MC0  MD  ME  OP4  OP3  OP2  OP1  OP0  LDMAHR1  LDMAHR0  LoadCNT  CCSP  CST  LDOHR  CLROHR  CR15-CR8  CR7-CR0


always @ (IN)

	case(IN)

		8'd0: OUT = 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd1: OUT = 64'b0000000011000000000100000001000000101000000000000000000000000000;
		8'd2: OUT = 64'b0000000011000000010001110001000000101000100000000000000000000000;
		8'd3: OUT = 64'b0000000101100000001001110000000000000000000000000000000000000011;
		8'd4: OUT = 64'b0000000100000001000000000000000000000000000000000000000000000001;
		8'd10: OUT = 64'b0000000010000000110000000000000011000000000000000000000000000001;
		8'd11: OUT = 64'b0000000010000000110000000000001011000000000000000000000000000001;
		8'd12: OUT = 64'b0000000010000000110000000100000011000000000000000000000000000001;
		8'd13: OUT = 64'b0000000010000000110000000100001011000000000000000000000000000001;
		8'd14: OUT = 64'b0000000010000000100000000000000011000000000000000000000000000001;
		8'd15: OUT = 64'b0000000010000000100000000000001011000000000000000000000000000001;
		8'd16: OUT = 64'b0000000011000000000100000000001000101010100000000000000000000000;
		8'd17: OUT = 64'b0000000101101011000001100000000000000000000000000001001000111111;
		8'd18: OUT = 64'b0000000101100000000011100000000000010000000000000000000000010010;
		8'd19: OUT = 64'b0000000010000000010000000000000011000000000000000000000000000001;
		8'd20: OUT = 64'b0000000010000000000100000000001000101011000000000000000000010001;
		/*0000000010000000000100000000000000101011100000000000000000010001
		0000000010000000000100000000001000101100000000000000000000010001
		0000000010000000010000000000001000101010100000000000000000010000
		0000000010000000010000000000001000101011000000000000000000010100
		0000000010000000010000000000000000101011100000000000000000010101
		0000000010000000010000000000000000101100000000000000000000010110
		0000000010000000000100000000000000000000000000000000000000100000
		0000000011000000000100000000000000000000000000000000000000000000
		0000000101101011000001100000000000000000000000000001111001000000
		0000000101100000000011100000000000010000000000000000000000011110
		0000000101010010010000000000000011000000000000000000000000110110
		0000000101101011000001100000000000000000000000000010000101000001
		0000000101100000000011100000000000010000000000000000000000100001
		0000000101010010010000000000000011000000000000000000000000111000
		0000000011000000000100000000001000101010100000000000000000000000
		0000000011000000000010000011000000000000000000000000000000000000
		0000000101101011000000100000000000000000000000000010011001000010
		0000000101101000000000100000000000000000000000000000000100100110
		0000000010000000000100000000001000101011000000000000000000100100
		0000000010000000000100000000000000101011100000000000000000100100
		0000000010000000000100000000000000101100000000000000000000100100
		0000000010000000010000000000001000101010100000000000000000100011
		0000000010000000010000000000001000101011000000000000000000100011
		0000000010000000010000000000000000101011100000000000000000101000
		0000000010000000010000000000000000101100000000000000000000101001
		0000000011000000000100000000000000101000000000000000000000000000
		0000000011000000000010000011000000000000000000000000000000000000
		0000000101101011000000100000000000000000000000000011000101000011
		0000000101101000000000100000000000000000000000000011100000110001
		0000000011000000000100000000000000101000000000000000000000000000
		0000000011000000000010000011000000000000000000000000000000000000
		0000000101101011000000100000000000000000000000000011010101000101
		0000000101101000000000100000000000000000000000000011011000110101
		0000000010000000010000000000000000101011100000000000000000000001
		0000000010000000010000000000000000101100000000000000000000000001
		0000000010000000010000000000001000101010100000000000000000000001
		0000000010000000010000000000001000101011000000000000000000000001
		0000000101101000000000100000000000000000000000000011100100111010
		0000000101101000000000100000000000000000000000000011011100111011
		0000000011000000000100000000000000101000000000000000000000000000
		0000000011000000000010000011000000000000000000000000000000000000
		0000000101101011000000100000000000000000000000000011101001000100
		0000000101101000000011110000000000010000000000000001001100111111
		0000000101101000000011110000000000010000000000000001111101000000
		0000000101101000000011110000000000010000000000000010001001000001
		0000000101101000000011110000000000010000000000000000000101000010
		0000000101101000000011110000000000010000000000000011100001000011
		0000000101101000000011110000000000010000000000000011100101000100
		0000000101101000000011110000000000010000000000000011011001000101
		0000000011000000000100000000000000101000000000000000000000000000
		0000000011000000000010000011000000000000000000000000000000000000
		0000000101101011000000100000000000000000000000000011101101001001
		0000000101101000000011110000000000010000000000000011011101001001
		0000000011000000000100001000001000101010100000000000000000000000
		0000000011000000000001101000000000000000000000000000000000000000
		0000000101100000000011101000000000010000000000000000000001001100
		0000000010000000010000001000000011000000000000000000000000000001
		0000000010000000000100001000001000101011000000000000000001001011
		0000000010000000000100001000000000101011100000000000000001001011
		0000000010000000000100001000001000101100000000000000000001001011
		0000000010000000010000001000001000101010100000000000000001001010
		0000000010000000010000001000001000101011000000000000000001001110
		0000000010000000010000001000000000101011100000000000000001001111
		0000000010000000010000001000000000101100000000000000000001010000
		0000000011000000000100001000000000000000000000000000000000000000
		0000000011000000000001101000000000000000000000000000000000000000
		0000000101100000000011101000000000010000000000000000000001010111
		0000000101100010010000001000000011000000000000000000000001011010
		0000000010000000010000001000000000101011100000000000000000000001
		0000000010000000010000001000000000101100000000000000000000000001
		0000000011000000000100001000000000000000000000000000000000000000
		0000000011000000000001101000000000000000000000000000000000000000
		0000000101100000000011101000000000010000000000000000000001011101
		0000000101100010010000001000000011000000000000000000000001100000
		0000000010000000010000001000001000101010100000000000000000000001
		0000000010000000010000001000001000101011000000000000000000000001
		0000000011000000000100001000001000101010100000000000000000000000
		0000000011000000000010001011000000000000000000000000000000000000
		0000000011000000000000101000000000000000000000000000000000000000
		0000000101101000000000101000000000000000000000000000000101100100
		0000000010000000000100001000001000101011000000000000000001100010
		0000000010000000000100001000000000101011100000000000000001100010
		0000000010000000000100001000000000101100000000000000000001100010
		0000000010000000010000001000001000101010100000000000000001100001
		0000000010000000010000001000001000101011000000000000000001100001
		0000000010000000010000001000000000101011100000000000000001100110
		0000000010000000010000001000000000101100000000000000000001100111
		0000000011000000000100001000000000101000000000000000000000000000
		0000000011000000000010001011000000000000000000000000000000000000
		0000000011000000000000101000000000000000000000000000000000000000
		0000000101101000000000101000000000000000000000000101111101101111
		0000000011000000000100001000000000101000000000000000000000000000
		0000000011000000000010001011000000000000000000000000000000000000
		0000000011000000000000101000000000000000000000000000000000000000
		0000000101101000000000101000000000000000000000000110000001110011
		0000000011000000000100001000000000101000000000000000000000000000
		0000000011000000000010001011000000000000000000000000000000000000
		0000000011000000000000101000000000000000000000000000000000000000
		0000000101101000000000101000000000000000000000000101100101110111
		0000000011000000000100001000000000101000000000000000000000000000
		0000000011000000000010001011000000000000000000000000000000000000
		0000000011000000000000101000000000000000000000000000000000000000
		0000000101101000000000101000000000000000000000000101101001111011
		0000000011000000000100011000001000101010100000000000000000000000
		0000000011000000000001111000000000000000000000000000000000000000
		0000000101100000000011111000000000010000000000000000000001111110
		0000000010000000010000011000000011000000000000000000000000000001
		0000000010000000000100011000001000101011000000000000000001111101
		0000000010000000000100011000000000101011100000000000000001111101
		0000000010000000000100011000001000101100000000000000000001111101
		0000000010000000010000011000001000101010100000000000000001111100
		0000000010000000010000011000001000101011000000000000000010000000
		0000000010000000010000011000000000101011100000000000000010000001
		0000000010000000010000011000000000101100000000000000000010000010
		0000000011000000000100011000000000000000000000000000000000000000
		0000000011000000000001111000000000000000000000000000000000000000
		0000000101100000000011111000000000010000000000000000000010001001
		0000000101100010010000011000000011000000000000000000000010001011
		0000000010000000010000011000000000101011100000000000000000000001
		0000000010000000010000011000000000101100000000000000000000000001
		0000000011000000000100011000000000000000000000000000000000000000
		0000000011000000000001111000000000000000000000000000000000000000
		0000000101100000000011111000000000010000000000000000000010001111
		0000000101100010010000011000000011000000000000000000000010010010
		0000000010000000010000011000001000101010100000000000000000000001
		0000000010000000010000011000001000101011000000000000000000000001
		0000000011000010000100011000001000101010100000000000000000000000
		0000000011000000000010011011000000000000000000000000000000000000
		0000000011000000000000111000000000000000000000000000000000000000
		0000000101101000000000111000000000000000000000000000000110010110
		0000000010000000000100011000001000101011000000000000000010010100
		0000000010000000000100011000000000101011100000000000000010010100
		0000000010000000000100011000000000101100000000000000000010010100
		0000000010000000010000011000001000101010100000000000000010010011
		0000000010000000010000011000001000101011000000000000000010010011
		0000000010000000010000011000000000101011100000000000000010011000
		0000000010000000010000011000000000101100000000000000000010011001
		0000000011000000000100011000000000101000000000000000000000000000
		0000000011000000000010011011000000000000000000000000000000000000
		0000000011000000000000111000000000000000000000000000000000000000
		0000000101101000000000111000000000000000000000001001000110100001
		0000000011000000000100011000000000101000000000000000000000000000
		0000000011000000000010011011000000000000000000000000000000000000
		0000000011000000000000111000000000000000000000000000000000000000
		0000000101101000000000111000000000000000000000001001001010100101
		0000000011000000000100011000000000101000000000000000000000000000
		0000000011000000000010011011000000000000000000000000000000000000
		0000000011000000000000111000000000000000000000000000000000000000
		0000000101101000000000111000000000000000000000001000101110101001
		0000000011000000000100011000000000101000000000000000000000000000
		0000000011000000000010011011000000000000000000000000000000000000
		0000000011000000000000111000000000000000000000000000000000000000
		0000000101101000000000111000000000000000000000001000110010101101
		0000000011000000000100011000001000101010100000000000000000000000
		0000000011000000000001111000000000000000000000000000000000000000
		0000000101100000000011111000000000010000000000000000000010110000
		0000000010000000010000011000000011000000000000000000000000000001
		0000000010000000000100011000001000101011000000000000000010101111
		0000000010000000000100011000000000101011100000000000000010101111
		0000000010000000000100011000001000101100000000000000000010101111
		0000000010000000010000011000001000101010100000000000000010101110
		0000000010000000010000011000001000101011000000000000000010110010
		0000000010000000010000011000000000101011100000000000000010110011
		0000000010000000010000011000000000101100000000000000000010110100
		0000000011000000000100011000000000000000000000000000000000000000
		0000000011000000000001111000000000000000000000000000000000000000
		0000000101100000000011111000000000010000000000000000000010111011
		0000000101100000010000011000000011000000000000000000000010111100
		0000000010000000010000011000000000101011100000000000000000000001
		0000000010000000010000011000000000101100000000000000000000000001
		0000000011000000000100011000000000000000000000000000000000000000
		0000000011000000000001111000000000000000000000000000000000000000
		0000000101100000000011111000000000010000000000000000000011000001
		0000000101100010010000011000000011000000000000000000000010111100
		0000000010000000010000011000001000101010100000000000000000000001
		0000000010000000010000011000001000101011000000000000000000000001
		0000000010000000000100000000000000101000111101010000000011001001
		0000000010000000000100000000000000101001011101010000000011001001
		0000000010000000000100000000000000101000111101010000000011001001
		0000000011000000000100000000000000101001011101010000000000000000
		0000000101100100000000000000000000000000010010100000000011010111
		0000000011000000000011110000000000110000000001000000000000000000
		0000000101100000010000000000010100101100100001000000000011001101
		0000000101101101000100000000010000101101000000011101011111001001
		0000000101101101000100000000010000101101100000011101011111001001
		0000000010000000000100000000000000101000111101010000000011010010
		0000000010000000000100000000000000101001011101010000000011010010
		0000000010000000000100000000000000101000111101010000000011010010
		0000000011000000000100000000000000101001011101010000000000000000
		0000000101100100000000000000000000000000010010100000000011010111
		0000000011000000000010000010000000101000000001000000000000000000
		0000000101100000000000110000000000000000000001000000000011010110
		0000000101101101000100000000010000101101000000011101011111010010
		0000000101101101000100000000010000101101100000011101011111010010
		0000000010000000010000000000011100101100100001000000000000000001
		0000000010000000010000000001001001101011100000000000000000000001
		0000000010000000010000000001000010101000000000000000000011011000
*/


	endcase //IN

endmodule //




//Duuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuureeeexxxxxxxxxxxxxxx!